module svm_ctrl #(
    parameter
) (
    input  [BID_W - 1 : 0] bid,
    
);
    
endmodule