module led_control #(
    parameters
) (
    port_list
);
    
endmodule