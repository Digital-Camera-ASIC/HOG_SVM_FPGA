package base_uvm_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "base_item.sv"
  `include "base_driver.sv"
  `include "base_monitor.sv"
  `include "base_agent.sv"
  `include "base_scoreboard.sv"
  `include "base_sequence.sv"
  `include "base_env.sv"
endpackage
